.source(Dark Web)
.search(bitcoin)
.find(.btc).column(btc addr)
.showRanges.showDate
.panel(Results)